module and_32bit(result,a,b);
input[31:0] a,b;
output [31:0] result;
	
and and0(result[0],a[0],b[0]);
and and1(result[1],a[1],b[1]);
and and2(result[2],a[2],b[2]);
and and3(result[3],a[3],b[3]);
and and4(result[4],a[4],b[4]);
and and5(result[5],a[5],b[5]);
and and6(result[6],a[6],b[6]);
and and7(result[7],a[7],b[7]);
and and8(result[8],a[8],b[8]);
and and9(result[9],a[9],b[9]);
and and10(result[10],a[10],b[10]);
and and11(result[11],a[11],b[11]);
and and12(result[12],a[12],b[12]);
and and13(result[13],a[13],b[13]);
and and14(result[14],a[14],b[14]);
and and15(result[15],a[15],b[15]);
and and16(result[16],a[16],b[16]);
and and17(result[17],a[17],b[17]);
and and18(result[18],a[18],b[18]);
and and19(result[19],a[19],b[19]);
and and20(result[20],a[20],b[20]);
and and21(result[21],a[21],b[21]);
and and22(result[22],a[22],b[22]);
and and23(result[23],a[23],b[23]);
and and24(result[24],a[24],b[24]);
and and25(result[25],a[25],b[25]);
and and26(result[26],a[26],b[26]);
and and27(result[27],a[27],b[27]);
and and28(result[28],a[28],b[28]);
and and29(result[29],a[29],b[29]);
and and30(result[30],a[30],b[30]);
and and31(result[31],a[31],b[31]);
	
endmodule